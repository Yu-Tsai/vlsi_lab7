//*************************************************                       
//** Author: LPHP Lab                               
//** Project: Simple image processor
//**    			- Grayscale
//*************************************************


module grayscale(clk,
                 rst,
                 en,
                 d,
                 q);

// ---------------------- input  ---------------------- //
  input clk;
  input rst;
  input en;
  input [23:0]d;
  
// ---------------------- output ---------------------- //  
  output reg[7:0]q;
// --------------- below is your design --------------- //
  

  
  
endmodule
// ------------------ the end of code ------------------ //